module score
  (
  curr_x,
  curr_y,
  key,


  );

  input [7:0] curr_x, curr_y;
  input [3:0] key;

  output [6:0] score;



  
